library ieee;
use ieee.std_logic_1164.all; -- use of std_logic

-- Next is the making of the entity.
entity full_adder_single_flip is
	port(
		-- Full adder inputs
		FA_a	: in std_logic;
		FA_b	: in std_logic;
		FA_cin	: in std_logic;
		-- Register necassary inputs
		clk		: in std_logic;
		rst_n	: in std_logic;
		-- space between inputs and outputs.
		-- Register outputs
		Reg_SumF	: out std_logic;
		Reg_coutF	: out std_logic
	);
end entity full_adder_single_flip;

architecture behave of full_adder_single_flip is
component full_adder is
	port( 
		a		: in std_logic; -- Full adder stuff.
		b		: in std_logic;
		cin		: in std_logic;
		-- space between inputs and outputs.
		sumF	: out std_logic;
		coutF	: out std_logic
		);
end component full_adder;

component d_flip_flop_signal is
	port( 
		Data 	: in std_logic;
		clk		: in std_logic;
		rst_n	: in std_logic;
		Q 		: out std_logic
		);
end component d_flip_flop_signal;

signal s1: std_logic; -- Intermediate signals for register and FA.
signal s2: std_logic; -- Intermediate signals

begin

-- cin has to be the and gate of a and x to work properly
FA: full_adder port map (
						a=>FA_a,
						b=>FA_b,
						cin=>FA_cin,
						sumF=>s1,
						coutF=>s2
						);
REG: d_flip_flop_signal port map (
						Data=>s1,
						clk=>clk,
						rst_n=>rst_n,
						Q=>Reg_SumF
						);
REG2: d_flip_flop_signal port map (
						Data=>s2,
						clk=>clk,
						rst_n=>rst_n,
						Q=>Reg_coutF
						);

end architecture behave;